//Verilog HDL for "COMP12111_lib", "quiz32" "functional"


module quiz32 (input	CLK, R, a,
	       output reg       s);
reg [1:0] next_st;


endmodule
